-- AESproject.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AESproject is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity AESproject;

architecture rtl of AESproject is
	component aes_accelerator is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			am_address     : out std_logic_vector(31 downto 0);                    -- address
			am_byteEnable  : out std_logic_vector(3 downto 0);                     -- byteenable
			am_write       : out std_logic;                                        -- write
			am_read        : out std_logic;                                        -- read
			am_writeData   : out std_logic_vector(31 downto 0);                    -- writedata
			am_readData    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			am_waitRequest : in  std_logic                     := 'X';             -- waitrequest
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			as_address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			as_chipSelect  : in  std_logic                     := 'X';             -- chipselect
			as_write       : in  std_logic                     := 'X';             -- write
			as_read        : in  std_logic                     := 'X';             -- read
			as_writeData   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			as_readData    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component aes_accelerator;

	component AESproject_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component AESproject_counter_0;

	component AESproject_epcs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic                                         -- irq
		);
	end component AESproject_epcs;

	component inv_aes_accelerator is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			as_address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			as_chipSelect  : in  std_logic                     := 'X';             -- chipselect
			as_write       : in  std_logic                     := 'X';             -- write
			as_read        : in  std_logic                     := 'X';             -- read
			as_writeData   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			as_readData    : out std_logic_vector(31 downto 0);                    -- readdata
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			am_address     : out std_logic_vector(31 downto 0);                    -- address
			am_byteEnable  : out std_logic_vector(3 downto 0);                     -- byteenable
			am_write       : out std_logic;                                        -- write
			am_read        : out std_logic;                                        -- read
			am_writeData   : out std_logic_vector(31 downto 0);                    -- writedata
			am_readData    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			am_waitRequest : in  std_logic                     := 'X'              -- waitrequest
		);
	end component inv_aes_accelerator;

	component AESproject_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component AESproject_jtag_uart_0;

	component AESproject_nios2_qsys_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component AESproject_nios2_qsys_0;

	component AESproject_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component AESproject_onchip_memory;

	component AESproject_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component AESproject_sysid_qsys_0;

	component AESproject_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component AESproject_timer_0;

	component AESproject_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                            : in  std_logic                     := 'X';             -- clk
			aes_accelerator_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			aes_accelerator_0_avalon_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			aes_accelerator_0_avalon_master_waitrequest              : out std_logic;                                        -- waitrequest
			aes_accelerator_0_avalon_master_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			aes_accelerator_0_avalon_master_read                     : in  std_logic                     := 'X';             -- read
			aes_accelerator_0_avalon_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			aes_accelerator_0_avalon_master_write                    : in  std_logic                     := 'X';             -- write
			aes_accelerator_0_avalon_master_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			inv_aes_accelerator_0_avalon_master_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			inv_aes_accelerator_0_avalon_master_waitrequest          : out std_logic;                                        -- waitrequest
			inv_aes_accelerator_0_avalon_master_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			inv_aes_accelerator_0_avalon_master_read                 : in  std_logic                     := 'X';             -- read
			inv_aes_accelerator_0_avalon_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			inv_aes_accelerator_0_avalon_master_write                : in  std_logic                     := 'X';             -- write
			inv_aes_accelerator_0_avalon_master_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_address                         : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest                     : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                            : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                           : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess                     : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address                  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest              : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read                     : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_instruction_master_readdatavalid            : out std_logic;                                        -- readdatavalid
			aes_accelerator_0_avalon_slave_address                   : out std_logic_vector(2 downto 0);                     -- address
			aes_accelerator_0_avalon_slave_write                     : out std_logic;                                        -- write
			aes_accelerator_0_avalon_slave_read                      : out std_logic;                                        -- read
			aes_accelerator_0_avalon_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			aes_accelerator_0_avalon_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			aes_accelerator_0_avalon_slave_chipselect                : out std_logic;                                        -- chipselect
			counter_0_control_slave_address                          : out std_logic_vector(2 downto 0);                     -- address
			counter_0_control_slave_write                            : out std_logic;                                        -- write
			counter_0_control_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			counter_0_control_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			counter_0_control_slave_begintransfer                    : out std_logic;                                        -- begintransfer
			epcs_epcs_control_port_address                           : out std_logic_vector(8 downto 0);                     -- address
			epcs_epcs_control_port_write                             : out std_logic;                                        -- write
			epcs_epcs_control_port_read                              : out std_logic;                                        -- read
			epcs_epcs_control_port_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			epcs_epcs_control_port_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			epcs_epcs_control_port_chipselect                        : out std_logic;                                        -- chipselect
			inv_aes_accelerator_0_avalon_slave_address               : out std_logic_vector(2 downto 0);                     -- address
			inv_aes_accelerator_0_avalon_slave_write                 : out std_logic;                                        -- write
			inv_aes_accelerator_0_avalon_slave_read                  : out std_logic;                                        -- read
			inv_aes_accelerator_0_avalon_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			inv_aes_accelerator_0_avalon_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			inv_aes_accelerator_0_avalon_slave_chipselect            : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                      : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                       : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                 : out std_logic;                                        -- chipselect
			nios2_qsys_0_debug_mem_slave_address                     : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_debug_mem_slave_write                       : out std_logic;                                        -- write
			nios2_qsys_0_debug_mem_slave_read                        : out std_logic;                                        -- read
			nios2_qsys_0_debug_mem_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_debug_mem_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_debug_mem_slave_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_debug_mem_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_debug_mem_slave_debugaccess                 : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                                 : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory_s1_write                                   : out std_logic;                                        -- write
			onchip_memory_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                                   : out std_logic;                                        -- clken
			sysid_qsys_0_control_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                         : out std_logic;                                        -- write
			timer_0_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                    : out std_logic;                                        -- chipselect
			timer_1_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                         : out std_logic;                                        -- write
			timer_1_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component AESproject_mm_interconnect_0;

	component AESproject_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component AESproject_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal aes_accelerator_0_avalon_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:aes_accelerator_0_avalon_master_readdata -> aes_accelerator_0:am_readData
	signal aes_accelerator_0_avalon_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:aes_accelerator_0_avalon_master_waitrequest -> aes_accelerator_0:am_waitRequest
	signal aes_accelerator_0_avalon_master_address                         : std_logic_vector(31 downto 0); -- aes_accelerator_0:am_address -> mm_interconnect_0:aes_accelerator_0_avalon_master_address
	signal aes_accelerator_0_avalon_master_byteenable                      : std_logic_vector(3 downto 0);  -- aes_accelerator_0:am_byteEnable -> mm_interconnect_0:aes_accelerator_0_avalon_master_byteenable
	signal aes_accelerator_0_avalon_master_read                            : std_logic;                     -- aes_accelerator_0:am_read -> mm_interconnect_0:aes_accelerator_0_avalon_master_read
	signal aes_accelerator_0_avalon_master_write                           : std_logic;                     -- aes_accelerator_0:am_write -> mm_interconnect_0:aes_accelerator_0_avalon_master_write
	signal aes_accelerator_0_avalon_master_writedata                       : std_logic_vector(31 downto 0); -- aes_accelerator_0:am_writeData -> mm_interconnect_0:aes_accelerator_0_avalon_master_writedata
	signal inv_aes_accelerator_0_avalon_master_readdata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:inv_aes_accelerator_0_avalon_master_readdata -> inv_aes_accelerator_0:am_readData
	signal inv_aes_accelerator_0_avalon_master_waitrequest                 : std_logic;                     -- mm_interconnect_0:inv_aes_accelerator_0_avalon_master_waitrequest -> inv_aes_accelerator_0:am_waitRequest
	signal inv_aes_accelerator_0_avalon_master_address                     : std_logic_vector(31 downto 0); -- inv_aes_accelerator_0:am_address -> mm_interconnect_0:inv_aes_accelerator_0_avalon_master_address
	signal inv_aes_accelerator_0_avalon_master_byteenable                  : std_logic_vector(3 downto 0);  -- inv_aes_accelerator_0:am_byteEnable -> mm_interconnect_0:inv_aes_accelerator_0_avalon_master_byteenable
	signal inv_aes_accelerator_0_avalon_master_read                        : std_logic;                     -- inv_aes_accelerator_0:am_read -> mm_interconnect_0:inv_aes_accelerator_0_avalon_master_read
	signal inv_aes_accelerator_0_avalon_master_write                       : std_logic;                     -- inv_aes_accelerator_0:am_write -> mm_interconnect_0:inv_aes_accelerator_0_avalon_master_write
	signal inv_aes_accelerator_0_avalon_master_writedata                   : std_logic_vector(31 downto 0); -- inv_aes_accelerator_0:am_writeData -> mm_interconnect_0:inv_aes_accelerator_0_avalon_master_writedata
	signal nios2_qsys_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_debugaccess                            : std_logic;                     -- nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_address                                : std_logic_vector(17 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_data_master_read                                   : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_write                                  : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                         : std_logic_vector(17 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                            : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal nios2_qsys_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	signal mm_interconnect_0_onchip_memory_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                     : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                      : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                        : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                        : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_chipselect     : std_logic;                     -- mm_interconnect_0:aes_accelerator_0_avalon_slave_chipselect -> aes_accelerator_0:as_chipSelect
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_readdata       : std_logic_vector(31 downto 0); -- aes_accelerator_0:as_readData -> mm_interconnect_0:aes_accelerator_0_avalon_slave_readdata
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:aes_accelerator_0_avalon_slave_address -> aes_accelerator_0:as_address
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_read           : std_logic;                     -- mm_interconnect_0:aes_accelerator_0_avalon_slave_read -> aes_accelerator_0:as_read
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_write          : std_logic;                     -- mm_interconnect_0:aes_accelerator_0_avalon_slave_write -> aes_accelerator_0:as_write
	signal mm_interconnect_0_aes_accelerator_0_avalon_slave_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:aes_accelerator_0_avalon_slave_writedata -> aes_accelerator_0:as_writeData
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_chipselect : std_logic;                     -- mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_chipselect -> inv_aes_accelerator_0:as_chipSelect
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_readdata   : std_logic_vector(31 downto 0); -- inv_aes_accelerator_0:as_readData -> mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_readdata
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_address    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_address -> inv_aes_accelerator_0:as_address
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_read       : std_logic;                     -- mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_read -> inv_aes_accelerator_0:as_read
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_write      : std_logic;                     -- mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_write -> inv_aes_accelerator_0:as_write
	signal mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:inv_aes_accelerator_0_avalon_slave_writedata -> inv_aes_accelerator_0:as_writeData
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	signal mm_interconnect_0_epcs_epcs_control_port_chipselect             : std_logic;                     -- mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	signal mm_interconnect_0_epcs_epcs_control_port_readdata               : std_logic_vector(31 downto 0); -- epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	signal mm_interconnect_0_epcs_epcs_control_port_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	signal mm_interconnect_0_epcs_epcs_control_port_read                   : std_logic;                     -- mm_interconnect_0:epcs_epcs_control_port_read -> mm_interconnect_0_epcs_epcs_control_port_read:in
	signal mm_interconnect_0_epcs_epcs_control_port_write                  : std_logic;                     -- mm_interconnect_0:epcs_epcs_control_port_write -> mm_interconnect_0_epcs_epcs_control_port_write:in
	signal mm_interconnect_0_epcs_epcs_control_port_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_counter_0_control_slave_readdata              : std_logic_vector(31 downto 0); -- counter_0:readdata -> mm_interconnect_0:counter_0_control_slave_readdata
	signal mm_interconnect_0_counter_0_control_slave_address               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:counter_0_control_slave_address -> counter_0:address
	signal mm_interconnect_0_counter_0_control_slave_begintransfer         : std_logic;                     -- mm_interconnect_0:counter_0_control_slave_begintransfer -> counter_0:begintransfer
	signal mm_interconnect_0_counter_0_control_slave_write                 : std_logic;                     -- mm_interconnect_0:counter_0_control_slave_write -> counter_0:write
	signal mm_interconnect_0_counter_0_control_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:counter_0_control_slave_writedata -> counter_0:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- epcs:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- timer_1:irq -> irq_mapper:receiver3_irq
	signal nios2_qsys_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:aes_accelerator_0_reset_sink_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [epcs:reset_req, nios2_qsys_0:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal nios2_qsys_0_debug_reset_request_reset                          : std_logic;                     -- nios2_qsys_0:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_epcs_epcs_control_port_read_ports_inv         : std_logic;                     -- mm_interconnect_0_epcs_epcs_control_port_read:inv -> epcs:read_n
	signal mm_interconnect_0_epcs_epcs_control_port_write_ports_inv        : std_logic;                     -- mm_interconnect_0_epcs_epcs_control_port_write:inv -> epcs:write_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [aes_accelerator_0:rst_n, counter_0:reset_n, epcs:reset_n, inv_aes_accelerator_0:rst_n, jtag_uart_0:rst_n, nios2_qsys_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, timer_1:reset_n]

begin

	aes_accelerator_0 : component aes_accelerator
		port map (
			clk            => clk_clk,                                                     --         clock.clk
			am_address     => aes_accelerator_0_avalon_master_address,                     -- avalon_master.address
			am_byteEnable  => aes_accelerator_0_avalon_master_byteenable,                  --              .byteenable
			am_write       => aes_accelerator_0_avalon_master_write,                       --              .write
			am_read        => aes_accelerator_0_avalon_master_read,                        --              .read
			am_writeData   => aes_accelerator_0_avalon_master_writedata,                   --              .writedata
			am_readData    => aes_accelerator_0_avalon_master_readdata,                    --              .readdata
			am_waitRequest => aes_accelerator_0_avalon_master_waitrequest,                 --              .waitrequest
			rst_n          => rst_controller_reset_out_reset_ports_inv,                    --    reset_sink.reset_n
			as_address     => mm_interconnect_0_aes_accelerator_0_avalon_slave_address,    --  avalon_slave.address
			as_chipSelect  => mm_interconnect_0_aes_accelerator_0_avalon_slave_chipselect, --              .chipselect
			as_write       => mm_interconnect_0_aes_accelerator_0_avalon_slave_write,      --              .write
			as_read        => mm_interconnect_0_aes_accelerator_0_avalon_slave_read,       --              .read
			as_writeData   => mm_interconnect_0_aes_accelerator_0_avalon_slave_writedata,  --              .writedata
			as_readData    => mm_interconnect_0_aes_accelerator_0_avalon_slave_readdata    --              .readdata
		);

	counter_0 : component AESproject_counter_0
		port map (
			clk           => clk_clk,                                                 --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			address       => mm_interconnect_0_counter_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_counter_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_counter_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_counter_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_counter_0_control_slave_writedata      --              .writedata
		);

	epcs : component AESproject_epcs
		port map (
			clk        => clk_clk,                                                  --               clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			reset_req  => rst_controller_reset_out_reset_req,                       --                  .reset_req
			address    => mm_interconnect_0_epcs_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_0_epcs_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_0_epcs_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_0_epcs_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_0_epcs_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_0_epcs_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_mapper_receiver2_irq                                  --               irq.irq
		);

	inv_aes_accelerator_0 : component inv_aes_accelerator
		port map (
			clk            => clk_clk,                                                         --         clock.clk
			as_address     => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_address,    --  avalon_slave.address
			as_chipSelect  => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_chipselect, --              .chipselect
			as_write       => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_write,      --              .write
			as_read        => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_read,       --              .read
			as_writeData   => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_writedata,  --              .writedata
			as_readData    => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_readdata,   --              .readdata
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --    reset_sink.reset_n
			am_address     => inv_aes_accelerator_0_avalon_master_address,                     -- avalon_master.address
			am_byteEnable  => inv_aes_accelerator_0_avalon_master_byteenable,                  --              .byteenable
			am_write       => inv_aes_accelerator_0_avalon_master_write,                       --              .write
			am_read        => inv_aes_accelerator_0_avalon_master_read,                        --              .read
			am_writeData   => inv_aes_accelerator_0_avalon_master_writedata,                   --              .writedata
			am_readData    => inv_aes_accelerator_0_avalon_master_readdata,                    --              .readdata
			am_waitRequest => inv_aes_accelerator_0_avalon_master_waitrequest                  --              .waitrequest
		);

	jtag_uart_0 : component AESproject_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	nios2_qsys_0 : component AESproject_nios2_qsys_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_qsys_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_qsys_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_qsys_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_qsys_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_qsys_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_qsys_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_qsys_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_qsys_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_qsys_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_qsys_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_qsys_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_qsys_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_qsys_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_qsys_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory : component AESproject_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	sysid_qsys_0 : component AESproject_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component AESproject_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                      --   irq.irq
		);

	timer_1 : component AESproject_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	mm_interconnect_0 : component AESproject_mm_interconnect_0
		port map (
			clk_0_clk_clk                                            => clk_clk,                                                         --                                          clk_0_clk.clk
			aes_accelerator_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                  -- aes_accelerator_0_reset_sink_reset_bridge_in_reset.reset
			aes_accelerator_0_avalon_master_address                  => aes_accelerator_0_avalon_master_address,                         --                    aes_accelerator_0_avalon_master.address
			aes_accelerator_0_avalon_master_waitrequest              => aes_accelerator_0_avalon_master_waitrequest,                     --                                                   .waitrequest
			aes_accelerator_0_avalon_master_byteenable               => aes_accelerator_0_avalon_master_byteenable,                      --                                                   .byteenable
			aes_accelerator_0_avalon_master_read                     => aes_accelerator_0_avalon_master_read,                            --                                                   .read
			aes_accelerator_0_avalon_master_readdata                 => aes_accelerator_0_avalon_master_readdata,                        --                                                   .readdata
			aes_accelerator_0_avalon_master_write                    => aes_accelerator_0_avalon_master_write,                           --                                                   .write
			aes_accelerator_0_avalon_master_writedata                => aes_accelerator_0_avalon_master_writedata,                       --                                                   .writedata
			inv_aes_accelerator_0_avalon_master_address              => inv_aes_accelerator_0_avalon_master_address,                     --                inv_aes_accelerator_0_avalon_master.address
			inv_aes_accelerator_0_avalon_master_waitrequest          => inv_aes_accelerator_0_avalon_master_waitrequest,                 --                                                   .waitrequest
			inv_aes_accelerator_0_avalon_master_byteenable           => inv_aes_accelerator_0_avalon_master_byteenable,                  --                                                   .byteenable
			inv_aes_accelerator_0_avalon_master_read                 => inv_aes_accelerator_0_avalon_master_read,                        --                                                   .read
			inv_aes_accelerator_0_avalon_master_readdata             => inv_aes_accelerator_0_avalon_master_readdata,                    --                                                   .readdata
			inv_aes_accelerator_0_avalon_master_write                => inv_aes_accelerator_0_avalon_master_write,                       --                                                   .write
			inv_aes_accelerator_0_avalon_master_writedata            => inv_aes_accelerator_0_avalon_master_writedata,                   --                                                   .writedata
			nios2_qsys_0_data_master_address                         => nios2_qsys_0_data_master_address,                                --                           nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest                     => nios2_qsys_0_data_master_waitrequest,                            --                                                   .waitrequest
			nios2_qsys_0_data_master_byteenable                      => nios2_qsys_0_data_master_byteenable,                             --                                                   .byteenable
			nios2_qsys_0_data_master_read                            => nios2_qsys_0_data_master_read,                                   --                                                   .read
			nios2_qsys_0_data_master_readdata                        => nios2_qsys_0_data_master_readdata,                               --                                                   .readdata
			nios2_qsys_0_data_master_write                           => nios2_qsys_0_data_master_write,                                  --                                                   .write
			nios2_qsys_0_data_master_writedata                       => nios2_qsys_0_data_master_writedata,                              --                                                   .writedata
			nios2_qsys_0_data_master_debugaccess                     => nios2_qsys_0_data_master_debugaccess,                            --                                                   .debugaccess
			nios2_qsys_0_instruction_master_address                  => nios2_qsys_0_instruction_master_address,                         --                    nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest              => nios2_qsys_0_instruction_master_waitrequest,                     --                                                   .waitrequest
			nios2_qsys_0_instruction_master_read                     => nios2_qsys_0_instruction_master_read,                            --                                                   .read
			nios2_qsys_0_instruction_master_readdata                 => nios2_qsys_0_instruction_master_readdata,                        --                                                   .readdata
			nios2_qsys_0_instruction_master_readdatavalid            => nios2_qsys_0_instruction_master_readdatavalid,                   --                                                   .readdatavalid
			aes_accelerator_0_avalon_slave_address                   => mm_interconnect_0_aes_accelerator_0_avalon_slave_address,        --                     aes_accelerator_0_avalon_slave.address
			aes_accelerator_0_avalon_slave_write                     => mm_interconnect_0_aes_accelerator_0_avalon_slave_write,          --                                                   .write
			aes_accelerator_0_avalon_slave_read                      => mm_interconnect_0_aes_accelerator_0_avalon_slave_read,           --                                                   .read
			aes_accelerator_0_avalon_slave_readdata                  => mm_interconnect_0_aes_accelerator_0_avalon_slave_readdata,       --                                                   .readdata
			aes_accelerator_0_avalon_slave_writedata                 => mm_interconnect_0_aes_accelerator_0_avalon_slave_writedata,      --                                                   .writedata
			aes_accelerator_0_avalon_slave_chipselect                => mm_interconnect_0_aes_accelerator_0_avalon_slave_chipselect,     --                                                   .chipselect
			counter_0_control_slave_address                          => mm_interconnect_0_counter_0_control_slave_address,               --                            counter_0_control_slave.address
			counter_0_control_slave_write                            => mm_interconnect_0_counter_0_control_slave_write,                 --                                                   .write
			counter_0_control_slave_readdata                         => mm_interconnect_0_counter_0_control_slave_readdata,              --                                                   .readdata
			counter_0_control_slave_writedata                        => mm_interconnect_0_counter_0_control_slave_writedata,             --                                                   .writedata
			counter_0_control_slave_begintransfer                    => mm_interconnect_0_counter_0_control_slave_begintransfer,         --                                                   .begintransfer
			epcs_epcs_control_port_address                           => mm_interconnect_0_epcs_epcs_control_port_address,                --                             epcs_epcs_control_port.address
			epcs_epcs_control_port_write                             => mm_interconnect_0_epcs_epcs_control_port_write,                  --                                                   .write
			epcs_epcs_control_port_read                              => mm_interconnect_0_epcs_epcs_control_port_read,                   --                                                   .read
			epcs_epcs_control_port_readdata                          => mm_interconnect_0_epcs_epcs_control_port_readdata,               --                                                   .readdata
			epcs_epcs_control_port_writedata                         => mm_interconnect_0_epcs_epcs_control_port_writedata,              --                                                   .writedata
			epcs_epcs_control_port_chipselect                        => mm_interconnect_0_epcs_epcs_control_port_chipselect,             --                                                   .chipselect
			inv_aes_accelerator_0_avalon_slave_address               => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_address,    --                 inv_aes_accelerator_0_avalon_slave.address
			inv_aes_accelerator_0_avalon_slave_write                 => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_write,      --                                                   .write
			inv_aes_accelerator_0_avalon_slave_read                  => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_read,       --                                                   .read
			inv_aes_accelerator_0_avalon_slave_readdata              => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_readdata,   --                                                   .readdata
			inv_aes_accelerator_0_avalon_slave_writedata             => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_writedata,  --                                                   .writedata
			inv_aes_accelerator_0_avalon_slave_chipselect            => mm_interconnect_0_inv_aes_accelerator_0_avalon_slave_chipselect, --                                                   .chipselect
			jtag_uart_0_avalon_jtag_slave_address                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,         --                      jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,           --                                                   .write
			jtag_uart_0_avalon_jtag_slave_read                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,            --                                                   .read
			jtag_uart_0_avalon_jtag_slave_readdata                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                                                   .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                                                   .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                                                   .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      --                                                   .chipselect
			nios2_qsys_0_debug_mem_slave_address                     => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address,          --                       nios2_qsys_0_debug_mem_slave.address
			nios2_qsys_0_debug_mem_slave_write                       => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write,            --                                                   .write
			nios2_qsys_0_debug_mem_slave_read                        => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read,             --                                                   .read
			nios2_qsys_0_debug_mem_slave_readdata                    => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata,         --                                                   .readdata
			nios2_qsys_0_debug_mem_slave_writedata                   => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata,        --                                                   .writedata
			nios2_qsys_0_debug_mem_slave_byteenable                  => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable,       --                                                   .byteenable
			nios2_qsys_0_debug_mem_slave_waitrequest                 => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest,      --                                                   .waitrequest
			nios2_qsys_0_debug_mem_slave_debugaccess                 => mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess,      --                                                   .debugaccess
			onchip_memory_s1_address                                 => mm_interconnect_0_onchip_memory_s1_address,                      --                                   onchip_memory_s1.address
			onchip_memory_s1_write                                   => mm_interconnect_0_onchip_memory_s1_write,                        --                                                   .write
			onchip_memory_s1_readdata                                => mm_interconnect_0_onchip_memory_s1_readdata,                     --                                                   .readdata
			onchip_memory_s1_writedata                               => mm_interconnect_0_onchip_memory_s1_writedata,                    --                                                   .writedata
			onchip_memory_s1_byteenable                              => mm_interconnect_0_onchip_memory_s1_byteenable,                   --                                                   .byteenable
			onchip_memory_s1_chipselect                              => mm_interconnect_0_onchip_memory_s1_chipselect,                   --                                                   .chipselect
			onchip_memory_s1_clken                                   => mm_interconnect_0_onchip_memory_s1_clken,                        --                                                   .clken
			sysid_qsys_0_control_slave_address                       => mm_interconnect_0_sysid_qsys_0_control_slave_address,            --                         sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                      => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,           --                                                   .readdata
			timer_0_s1_address                                       => mm_interconnect_0_timer_0_s1_address,                            --                                         timer_0_s1.address
			timer_0_s1_write                                         => mm_interconnect_0_timer_0_s1_write,                              --                                                   .write
			timer_0_s1_readdata                                      => mm_interconnect_0_timer_0_s1_readdata,                           --                                                   .readdata
			timer_0_s1_writedata                                     => mm_interconnect_0_timer_0_s1_writedata,                          --                                                   .writedata
			timer_0_s1_chipselect                                    => mm_interconnect_0_timer_0_s1_chipselect,                         --                                                   .chipselect
			timer_1_s1_address                                       => mm_interconnect_0_timer_1_s1_address,                            --                                         timer_1_s1.address
			timer_1_s1_write                                         => mm_interconnect_0_timer_1_s1_write,                              --                                                   .write
			timer_1_s1_readdata                                      => mm_interconnect_0_timer_1_s1_readdata,                           --                                                   .readdata
			timer_1_s1_writedata                                     => mm_interconnect_0_timer_1_s1_writedata,                          --                                                   .writedata
			timer_1_s1_chipselect                                    => mm_interconnect_0_timer_1_s1_chipselect                          --                                                   .chipselect
		);

	irq_mapper : component AESproject_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_qsys_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_qsys_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_epcs_epcs_control_port_read_ports_inv <= not mm_interconnect_0_epcs_epcs_control_port_read;

	mm_interconnect_0_epcs_epcs_control_port_write_ports_inv <= not mm_interconnect_0_epcs_epcs_control_port_write;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of AESproject
